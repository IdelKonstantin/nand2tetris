/**
 * The ALU (Arithmetic Logic Unit).
 * Computes one of the following functions:
 * x+y, x-y, y-x, 0, 1, -1, x, y, -x, -y, !x, !y,
 * x+1, y+1, x-1, y-1, x&y, x|y on two 16-bit inputs,
 * according to 6 input bits denoted zx,nx,zy,ny,f,no.
 * In addition, the ALU computes two 1-bit outputs:
 * if the ALU output == 0, zr is set to 1; otherwise zr is set to 0;
 * if the ALU output < 0, ng is set to 1; otherwise ng is set to 0.
 */

// Implementation: the ALU logic manipulates the x and y inputs
// and operates on the resulting values, as follows:
// if (zx == 1) set x = 0        // 16-bit constant
// if (nx == 1) set x = !x       // bitwise not
// if (zy == 1) set y = 0        // 16-bit constant
// if (ny == 1) set y = !y       // bitwise not
// if (f == 1)  set out = x + y  // integer 2's complement addition
// if (f == 0)  set out = x & y  // bitwise and
// if (no == 1) set out = !out   // bitwise not
// if (out == 0) set zr = 1
// if (out < 0) set ng = 1

//`include "../mux2in1_16/mux2in1_16.v"

module ALU 
(
	input [15:0] x,
	input [15:0] y,
	input zx, zy, nx, ny, f, no,
	output [15:0] out,
	output zr,
	output ng
);

wire [15:0] zxMuxOut, zyMuxOut;
wire [15:0] notZxMuxOut, notZyMuxOut;
wire [15:0] nxMuxOut, nyMuxOut;
wire [15:0] addOut, andOut;
wire [15:0] fMuxOut, noFMuxOut;

wire highOr, lowOr;

mux2in1_16 zxMux(.a(x), .b(16'b0), .sel(zx), .y(zxMuxOut));
not_16 notzxMux(.a(zxMuxOut), .y(notZxMuxOut));
mux2in1_16 nxMux(.a(zxMuxOut), .b(notZxMuxOut), .sel(nx), .y(nxMuxOut));

mux2in1_16 zyMux(.a(y), .b(16'b0), .sel(zy), .y(zyMuxOut));
not_16 notZyMux(.a(zyMuxOut), .y(notZyMuxOut));
mux2in1_16 nyMux(.a(zyMuxOut), .b(notZyMuxOut), .sel(ny), .y(nyMuxOut));

add_16 assNxNy(.a(nxMuxOut), .b(nyMuxOut), .y(addOut));
and_16 andNxNy(.a(nxMuxOut), .b(nyMuxOut), .y(andOut));

mux2in1_16 fMux(.a(andOut), .b(addOut), .sel(f), .y(fMuxOut));
not_16 notFMux(.a(fMuxOut), .y(noFMuxOut));

mux2in1_16 noMux(.a(fMuxOut), .b(noFMuxOut), .sel(no), .y(out));

assign ng = out[15];

or8in1 orHighBits(.a(out[7:0]), .y(highOr));
or8in1 orLowBits(.a(out[15:8]), .y(lowOr));

assign anyBitsTrue = highOr | lowOr;
assign zr = ~anyBitsTrue;

endmodule